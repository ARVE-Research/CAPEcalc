netcdf MERRA2-CAPE {
dimensions:
	time = UNLIMITED ;
	lon = 576 ;
	lat = 361 ;
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1980-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	short CAPE(time, lat, lon) ;
		CAPE:long_name = "Convective Available Potential Energy" ;
		CAPE:units = "J kg-1" ;
		CAPE:_FillValue = -32768s ;
		CAPE:missing_value = -32768s ;
		CAPE:actual_range = 9999.f, -9999.f ;
		CAPE:scale_factor = 0.1f ;
		CAPE:add_offset = 3276.7f ;
		CAPE:_Storage = "chunked" ;
		CAPE:_ChunkSizes = 1, 361, 576 ;
		CAPE:_Shuffle = "true" ;
		CAPE:_DeflateLevel = 1 ;
	short CIN(time, lat, lon) ;
		CIN:long_name = "Convective Inhibition" ;
		CIN:units = "J kg-1" ;
		CIN:_FillValue = -32768s ;
		CIN:missing_value = -32768s ;
		CIN:actual_range = 9999.f, -9999.f ;
		CIN:scale_factor = 0.1f ;
		CIN:add_offset = 3276.7f ;
		CIN:_Storage = "chunked" ;
		CIN:_ChunkSizes = 1, 361, 576 ;
		CIN:_Shuffle = "true" ;
		CIN:_DeflateLevel = 1 ;

// global attributes:
		:Conventions = "COARDS, CF-1.11" ;
		:title = "MERRA2 estimated CAPE and CIN" ;
		:note = "calculated with NCAR getcape.f90" ;
		:node_offset = 1 ;
}
